verilog module
git